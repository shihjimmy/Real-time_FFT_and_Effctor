module Wrapper (
    input          avm_rst,
    input          avm_clk,
    output [  4:0] avm_address,
    output         avm_read,
    input  [ 31:0] avm_readdata,
    output         avm_write,
    output [ 31:0] avm_writedata,
    input          avm_waitrequest,
    // frequencies to sent
    input  [255:0] freqs,            // 16 16bit frequency amplitude 
    input          fft_ready,
    // parameters
    output [ 15:0] threshold_gate,   // -inf ~ 0 (0 ~ 32767)
    output [ 15:0] threshold_comp,   // -inf ~ 0 (0 ~ 32767)
    output [  4:0] ratio,            // 1:1 ~ 31:1
    output [ 15:0] makeup,           // (0 ~ 32767)
    output         GetMusic,
    output [  2:0] Pan
);

  localparam RX_BASE = 0 * 4;
  localparam TX_BASE = 1 * 4;
  localparam STATUS_BASE = 2 * 4;
  localparam TX_OK_BIT = 6;
  localparam RX_OK_BIT = 7;

  // States
  localparam S_IDLE = 0;
  localparam S_RECEIVE = 1;
  localparam S_SEND = 2;
  localparam S_UPDATE = 3;

  // parameters and frequencies
  logic [255:0] freqs_r, freqs_w;
  logic [15:0] threshold_gate_r, threshold_gate_w;
  logic [15:0] threshold_camp_r, threshold_camp_w;
  logic [4:0] ratio_r, ratio_w;
  logic [15:0] makeup_r, makeup_w;
  logic [2:0]  Pan_r, Pan_w;
  logic get_r, get_w;

  logic [1:0] state_r, state_w;
  logic [31:0] rcv_data_r, rcv_data_w;  // [31:16] id + [15:0] data
  logic [1:0] rcv_counter_r, rcv_counter_w;  // at most 4 bytes
  logic [4:0] send_counter_r, send_counter_w;  // at most 32 bytes
  logic [4:0] avm_address_r, avm_address_w;
  logic avm_read_r, avm_read_w, avm_write_r, avm_write_w;

  assign threshold_comp = threshold_camp_r;
  assign threshold_gate = threshold_gate_r;
  assign ratio = ratio_r;
  assign makeup = makeup_r;
  assign GetMusic = get_r;
  assign Pan = Pan_r;

  assign avm_address = avm_address_r;
  assign avm_read = avm_read_r;
  assign avm_write = avm_write_r;
  assign avm_writedata = freqs_r[255-:8];

  task StartRead;
    input [4:0] addr;
    begin
      avm_read_w = 1;
      avm_write_w = 0;
      avm_address_w = addr;
    end
  endtask

  task StartWrite;
    input [4:0] addr;
    begin
      avm_read_w = 0;
      avm_write_w = 1;
      avm_address_w = addr;
    end
  endtask

  always_comb begin
    get_w = 0;
    state_w = state_r;
    rcv_counter_w = rcv_counter_r;
    send_counter_w = send_counter_r;
    rcv_data_w = rcv_data_r;
    avm_address_w = avm_address_r;
    avm_read_w = avm_read_r;
    avm_write_w = avm_write_r;
    state_w = state_r;
    rcv_counter_w = rcv_counter_r;
    send_counter_w = send_counter_r;

    // parameters and frequencies
    freqs_w = freqs_r;
    threshold_gate_w = threshold_gate_r;
    threshold_camp_w = threshold_camp_r;
    ratio_w = ratio_r;
    makeup_w = makeup_r;
    Pan_w = Pan_r;

    case (state_r)
      S_IDLE: begin
        if (!avm_waitrequest && avm_readdata[RX_OK_BIT] && avm_address == STATUS_BASE) begin  // Rx ready => python ready to write
          state_w = S_RECEIVE;
          send_counter_w = 0;
          StartRead(RX_BASE);
        end 
        else if (!avm_waitrequest && avm_readdata[TX_OK_BIT] && avm_address == STATUS_BASE) begin  // Tx ready => python ready to read
          if (fft_ready) begin
            state_w = S_SEND;
            //when counter==0 loads frequency generated by FFT
            if (send_counter_r == 0) begin
              freqs_w = freqs;
            end
            StartWrite(TX_BASE);
          end
        end
        else begin
          // Rx isn't ready, do nothing
          state_w = S_IDLE;
        end
      end

      S_RECEIVE: begin
        if (!avm_waitrequest && avm_address == RX_BASE) begin
          StartRead(STATUS_BASE);
          rcv_data_w = (rcv_data_r << 8) + avm_readdata[7:0];
          if (&rcv_counter_r) begin  // finished
            state_w = S_UPDATE;
            rcv_counter_w = 2'd0;
          end 
          else begin
            state_w = S_IDLE;
            rcv_counter_w = rcv_counter_r + 2'd1;
          end
        end 
        else begin
          state_w = S_RECEIVE;
        end
      end

      S_SEND: begin
        if (!avm_waitrequest && avm_address == TX_BASE) begin
          StartRead(STATUS_BASE);
          freqs_w = freqs_r << 8;
          state_w = S_IDLE;
          if (&send_counter_r) begin  // finished
            send_counter_w = 0;
          end 
          else begin
            send_counter_w = send_counter_r + 5'd1;
          end
        end 
        else begin
          state_w = S_SEND;
        end
      end

      S_UPDATE: begin
        state_w = S_IDLE;

        rcv_data_w = rcv_data_r;
        StartRead(STATUS_BASE);
        case (rcv_data_r[31:16])
          16'd0: begin  // threshold (gate)
            threshold_gate_w = rcv_data_r[14:0];
          end
          16'd1: begin  // threshold (compressor)
            threshold_camp_w = rcv_data_r[14:0];
          end
          16'd2: begin  // ratio
            ratio_w = rcv_data_r[4:0];
          end
          16'd3: begin  // makeup
            makeup_w = rcv_data_r[14:0];
          end
          16'd4: begin
            Pan_w = rcv_data_r[2:0];
          end
          default: begin
            get_w = 1;
          end
        endcase
      end

    endcase
  end

  always_ff @(posedge avm_clk or posedge avm_rst) begin
    if (avm_rst) begin  // reset
      get_r <= 0;
      avm_address_r <= STATUS_BASE;
      avm_read_r <= 1;
      avm_write_r <= 0;
      state_r <= S_IDLE;
      rcv_counter_r <= 0;
      send_counter_r <= 0;
      rcv_data_r <= 32'd0;

      // parameters and frequencies
      freqs_r <= 0;
      makeup_r <= 1;
      threshold_gate_r <= 15'd1;
      threshold_camp_r <= 15'd16383;
      ratio_r <= 5;
      Pan_r <= 2;
    end 
    else begin
      get_r <= get_w;
      avm_address_r <= avm_address_w;
      avm_read_r <= avm_read_w;
      avm_write_r <= avm_write_w;
      state_r <= state_w;
      rcv_counter_r <= rcv_counter_w;
      send_counter_r <= send_counter_w;
      rcv_data_r <= rcv_data_w;

      // parameters and frequencies
      freqs_r <= freqs_w;
      makeup_r <= makeup_w;
      threshold_gate_r <= threshold_gate_w;
      threshold_camp_r <= threshold_camp_w;
      ratio_r <= ratio_w;
      Pan_r <= Pan_w;
    end
  end

endmodule